`define HADDR_SIZE 8 
`define HDATA_SIZE 32
